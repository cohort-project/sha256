package sha256_pkg;
    localparam  SHA_IF_DATA_W = 256;
    localparam  SHA256_DIGEST_W = 256;
    localparam  SHA256_BLOCK_W = 512;

endpackage