`ifndef SHA256_DEFS_SVH
`define SHA256_DEFS_SVH
    import sha256_pkg::*;
`endif